`timescale 1ns/1ps

module uart_irq_code_tb();

sim_top u_sim_top();

always begin
    if (
        u_sim_top.w_cpu_addr == 16'h0 &&
        u_sim_top.w_cpu_we == '1
    ) begin
        if (u_sim_top.w_cpu_data_from_cpu == 8'h6d) begin
            $display("Good finish!");
            $finish();
        end else begin
            $display("Bad finish!");
            $finish_and_return(-1);
        end
    end
    # 1;
end

initial begin
    repeat(15000) @(posedge u_sim_top.r_clk_cpu)
    u_sim_top.u_sim_uart.tx_en = 1;
    @(posedge u_sim_top.r_clk_cpu);
    u_sim_top.u_sim_uart.tx_data = 8'hAA;
    repeat (100) @(posedge u_sim_top.r_clk_cpu);
    $finish();
end

always @(u_sim_top.u_dut.u_rtc.r_output) begin
    $display("counter: %d", u_sim_top.u_dut.u_rtc.r_output);
end

endmodule