module sim_top();

//TODO: this
cpu_65c02 u_cpu();

//TODO: also this
super6502 u_dut();

//TODO: decide what to do here
memory u_mem();

endmodule