
localparam fSYS_MHz = 100;
localparam fCK_MHz  = 200;
localparam tIORT_u = 2;
localparam BL = 1;
localparam DDIO_TYPE = "SOFT";
localparam DQ_WIDTH  = 8;
localparam DQ_GROUP = 4;
localparam BA_WIDTH  = 2;
localparam ROW_WIDTH  = 13;
localparam COL_WIDTH  = 10;
localparam tPWRUP  = 200000;
localparam tRAS  = 44;
localparam tRC  = 66;
localparam tRCD = 20;
localparam tREF  = 64000000;
localparam tWR = 2;
localparam tMRD = 2;
localparam tRFC  = 66;
localparam tRAS_MAX = 120000;
localparam DATA_RATE = 2;
localparam tRP = 20;
localparam CL = 3;
