module sdram_adapter(
    input   i_sysclk,
    input   i_sdrclk,
    input   i_tACclk,
    input   i_pll_locked,
    output  o_pll_reset,
    output  o_sdr_CKE,
    output  o_sdr_n_CS,
    output  o_sdr_n_WE,
    output  o_sdr_n_RAS,
    output  o_sdr_n_CAS,
    output  [1:0]o_sdr_BA,
    output  [12:0]o_sdr_ADDR,
    input   [15:0]i_sdr_DATA,
    output  [15:0]o_sdr_DATA,
    output  [15:0]o_sdr_DATA_oe,
    output  [1:0]o_sdr_DQM
);

sdram u_sdram (
    .i_arst             (w_areset),
    .i_sysclk           (w_sysclk),
    .i_sdrclk           (i_sdrclk),
    .i_tACclk           (i_tACclk),
    .i_pll_locked       (1'b1),

    .i_we               (r_we_1P),
    .i_re               (r_re_1P),
    .i_last             (r_last_1P),
    .i_addr             (r_addr_1P),
    .i_din              (r_din_1P),
    .o_dout             (w_dout),
    .o_sdr_state        (w_sdr_state),
    .o_sdr_init_done    (w_sdr_init_done),
    .o_wr_ack           (w_wr_ack),
    .o_rd_ack           (w_rd_ack),
    .o_ref_req          (),
    .o_rd_valid         (w_rd_valid),

    .o_sdr_CKE          (w_sdr_CKE),
    .o_sdr_n_CS         (w_sdr_n_CS),
    .o_sdr_n_RAS        (w_sdr_n_RAS),
    .o_sdr_n_CAS        (w_sdr_n_CAS),
    .o_sdr_n_WE         (w_sdr_n_WE),
    .o_sdr_BA           (w_sdr_BA),
    .o_sdr_ADDR         (w_sdr_ADDR),
    .o_sdr_DATA         (w_sdr_DATA),
    .o_sdr_DATA_oe      (w_sdr_DATA_oe),
    .i_sdr_DATA         ({{16{1'b0}}, i_sdr_DATA}),
    .o_sdr_DQM          (w_sdr_DQM),

    .o_dbg_dly_cnt_b    (w_dbg_dly_cnt_b),
    .o_dbg_tRCD_done    (w_dbg_tRCD_done),
    .o_dbg_tRTW_done    (w_dbg_tRTW_done),
    .o_dbg_ref_req      (w_dbg_ref_req),
    .o_dbg_wr_ack       (w_dbg_wr_ack),
    .o_dbg_rd_ack       (w_dbg_rd_ack),
    .o_dbg_n_CS         (w_dbg_n_CS),
    .o_dbg_n_RAS        (w_dbg_n_RAS),
    .o_dbg_n_CAS        (w_dbg_n_CAS),
    .o_dbg_n_WE         (w_dbg_n_WE),
    .o_dbg_BA           (w_dbg_BA),
    .o_dbg_ADDR         (w_dbg_ADDR),
    .o_dbg_DATA_out     (w_dbg_DATA_out),
    .o_dbg_DATA_in      (w_dbg_DATA_in)
);

endmodule
